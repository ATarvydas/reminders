module buffer(
              input  A,
              output B);

   assign B = A;
   
   
endmodule
